// Copyright (c) 2017 Connectal Project

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

interface FastEchoIndication;
    method Action indication(Bit#(64) x);
endinterface

interface FastEchoRequest;
    method Action request(Bit#(64) x);
endinterface

interface FastEcho;
   interface FastEchoRequest request;
endinterface

module mkFastEcho#(FastEchoIndication indication)(FastEcho);
    Reg#(Maybe#(Bit#(64))) reqReg <- mkReg(tagged Invalid);

    rule sendIndication(reqReg matches tagged Valid .x);
        indication.indication(x);
        reqReg <= tagged Invalid;
    endrule

    interface FastEchoRequest request;
        method Action request(Bit#(64) x) if (!isValid(reqReg));
            reqReg <= tagged Valid x;
        endmethod
    endinterface
endmodule
